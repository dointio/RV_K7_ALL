module clk_wiz_0
   (clk_out1,
    clk_out2,
    clk_out3,
    resetn,
    locked,
    clk_in1);
  output clk_out1;
  output clk_out2;
  output clk_out3;
  input resetn;
  output locked;
  input clk_in1;

endmodule
